module ysyx_23060187_WBU(
    
);

endmodule