module numdisplay(
        input [31:0] num1,
        input [31:0] num2,
        input [31:0] num3,
        input [31:0] num4,
        input [31:0] num5,
        input [31:0] num6,
        input [31:0] num7,
        input [31:0] num8,
        output reg [6:0] seg1,
        output reg [6:0] seg2,
        output reg [6:0] seg3,
        output reg [6:0] seg4,
        output reg [6:0] seg5,
        output reg [6:0] seg6,
        output reg [6:0] seg7,
        output reg [6:0] seg8
    );

    always @(*) begin
        case(num1)
            32'h00000000:
                seg1 = 7'b0000001;
            32'h00000001:
                seg1 = 7'b1001111;
            32'h00000002:
                seg1 = 7'b0010010;
            32'h00000003:
                seg1 = 7'b0000110;
            32'h00000004:
                seg1 = 7'b1001100;
            32'h00000005:
                seg1 = 7'b0100100;
            32'h00000006:
                seg1 = 7'b0100000;
            32'h00000007:
                seg1 = 7'b0001111;
            32'h00000008:
                seg1 = 7'b0000000;
            32'h00000009:
                seg1 = 7'b0000100;
            default:
                seg1 = 7'b1111111;
        endcase
        case(num2)
            32'h00000000:
                seg2 = 7'b0000001;
            32'h00000001:
                seg2 = 7'b1001111;
            32'h00000002:
                seg2 = 7'b0010010;
            32'h00000003:
                seg2 = 7'b0000110;
            32'h00000004:
                seg2 = 7'b1001100;
            32'h00000005:
                seg2 = 7'b0100100;
            32'h00000006:
                seg2 = 7'b0100000;
            32'h00000007:
                seg2 = 7'b0001111;
            32'h00000008:
                seg2 = 7'b0000000;
            32'h00000009:
                seg2 = 7'b0000100;
            default:
                seg2 = 7'b1111111;
        endcase
        case(num3)
            32'h00000000:
                seg3 = 7'b0000001;
            32'h00000001:
                seg3 = 7'b1001111;
            32'h00000002:
                seg3 = 7'b0010010;
            32'h00000003:
                seg3 = 7'b0000110;
            32'h00000004:
                seg3 = 7'b1001100;
            32'h00000005:
                seg3 = 7'b0100100;
            32'h00000006:
                seg3 = 7'b0100000;
            32'h00000007:
                seg3 = 7'b0001111;
            32'h00000008:
                seg3 = 7'b0000000;
            32'h00000009:
                seg3 = 7'b0000100;
            default:
                seg3 = 7'b1111111;
        endcase
        case(num4)
            32'h00000000:
                seg4 = 7'b0000001;
            32'h00000001:
                seg4 = 7'b1001111;
            32'h00000002:
                seg4 = 7'b0010010;
            32'h00000003:
                seg4 = 7'b0000110;
            32'h00000004:
                seg4 = 7'b1001100;
            32'h00000005:
                seg4 = 7'b0100100;
            32'h00000006:
                seg4 = 7'b0100000;
            32'h00000007:
                seg4 = 7'b0001111;
            32'h00000008:
                seg4 = 7'b0000000;
            32'h00000009:
                seg4 = 7'b0000100;
            default:
                seg4 = 7'b1111111;
        endcase
        case(num5)
            32'h00000000:
                seg5 = 7'b0000001;
            32'h00000001:
                seg5 = 7'b1001111;
            32'h00000002:
                seg5 = 7'b0010010;
            32'h00000003:
                seg5 = 7'b0000110;
            32'h00000004:
                seg5 = 7'b1001100;
            32'h00000005:
                seg5 = 7'b0100100;
            32'h00000006:
                seg5 = 7'b0100000;
            32'h00000007:
                seg5 = 7'b0001111;
            32'h00000008:
                seg5 = 7'b0000000;
            32'h00000009:
                seg5 = 7'b0000100;
            default:
                seg5 = 7'b1111111;
        endcase
        case(num6)
            32'h00000000:
                seg6 = 7'b0000001;
            32'h00000001:
                seg6 = 7'b1001111;
            32'h00000002:
                seg6 = 7'b0010010;
            32'h00000003:
                seg6 = 7'b0000110;
            32'h00000004:
                seg6 = 7'b1001100;
            32'h00000005:
                seg6 = 7'b0100100;
            32'h00000006:
                seg6 = 7'b0100000;
            32'h00000007:
                seg6 = 7'b0001111;
            32'h00000008:
                seg6 = 7'b0000000;
            32'h00000009:
                seg6 = 7'b0000100;
            default:
                seg6 = 7'b1111111;
        endcase
        case(num7)
            32'h00000000:
                seg7 = 7'b0000001;
            32'h00000001:
                seg7 = 7'b1001111;
            32'h00000002:
                seg7 = 7'b0010010;
            32'h00000003:
                seg7 = 7'b0000110;
            32'h00000004:
                seg7 = 7'b1001100;
            32'h00000005:
                seg7 = 7'b0100100;
            32'h00000006:
                seg7 = 7'b0100000;
            32'h00000007:
                seg7 = 7'b0001111;
            32'h00000008:
                seg7 = 7'b0000000;
            32'h00000009:
                seg7 = 7'b0000100;
            default:
                seg7 = 7'b1111111;
        endcase
        case(num8)
            32'h00000000:
                seg8 = 7'b0000001;
            32'h00000001:
                seg8 = 7'b1001111;
            32'h00000002:
                seg8 = 7'b0010010;
            32'h00000003:
                seg8 = 7'b0000110;
            32'h00000004:
                seg8 = 7'b1001100;
            32'h00000005:
                seg8 = 7'b0100100;
            32'h00000006:
                seg8 = 7'b0100000;
            32'h00000007:
                seg8 = 7'b0001111;
            32'h00000008:
                seg8 = 7'b0000000;
            32'h00000009:
                seg8 = 7'b0000100;
            default:
                seg8 = 7'b1111111;
        endcase
    end

endmodule
